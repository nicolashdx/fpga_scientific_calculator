-- keyboard file