-- main file