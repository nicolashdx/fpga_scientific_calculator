-- alu file